// FIle Name:	lab2.sv
// Description:	Main for BCIT ELEX 7660, Lab 2.
//				This main file and its modules
//				Monitor for a keypress on a 4x4
//				keypad and then output the correct
//				keypress value to an LED screen
// Author:	Neil deHoog
// Date:		2018-01-19

module fish ( output logic [3:0] kpc,	// column select, active-low
			(* altera_attribute = "-name WEAK_PULL_UP_RESISTOR ON" *)
            input logic  [3:0] kpr, 	// rows, active-low w/ pull-ups
            output logic [7:0] leds,	// active-low LED segments 
            output logic [3:0] ct,  	// " digit enables
				output logic toggle_in,		// Input to the toggle switch. Always High
				input logic toggle_out, 	// Output from the toggle switch. Requires a pull up or down resistor
            input logic reset_n, CLOCK_50,
				output logic proximity_in,
				input logic proximity_out,
				output logic LED1,
				output logic LED2,
				output logic LED3,
				output logic LED4,
				output logic LED5,
				output logic LED6,
				output logic LED7,
				output logic LED8,
				output logic line_a,
				output logic line_b,
				output logic line_c,
				output logic line_d,
				input logic PW,
				output logic trig,
				input logic echo);

	logic clk ;                // 2kHz clock for keypad scanning
	logic kphit ;              // a key is pressed
	logic [3:0] num ;     		// value of pressed key
	logic [3:0] num_const = 0;	// stored value of the last pressed key
	logic toggle;					// logic value of the output from the toggle switch
	logic proximity;				// logic value of the input from the proximity sensor
	logic [1:0] dir = 2'b00;	// Motor direction variable
	logic [3:0] signal;			// Motor driver control signal
	logic [39:0] distance;
	logic [31:0] dist_test;
	logic [31:0] leng_test;
		
	
	assign ct = { {3{1'b0}}, 1'b1 } ;
	assign toggle_in = 0;
	assign proximity_in = 1;
   
	pll pll0 ( .inclk0(CLOCK_50), .c0(clk) ) ;
	decode7	decode7_0	(.num_const, .leds);
	kpdecode	kpdecode_0	(.kpc, .kpr, .kphit, .num, .num_const, .clk, .reset_n);
	colseq	colseq_0	(.kpr, .clk, .reset_n, .kpc);
	mode mode_0	(.toggle_out, .toggle, .clk, .LED1);
	optics optics_0 (.LED2, .proximity_out, .proximity, .clk);
	motor motor_0 (.clk, .reset_n, .dir, .signal);
	motor_decode motor_decode_0 (.signal, .clk, .line_a, .line_b, .line_c, .line_d);
	control control_0 (.clk, .toggle, .reset_n, .num, .num_const, .distance, .dir, .proximity_out, .dist_test, .leng_test);
	pulse pulse_0 (.clk, .trig, .echo, .distance);
		
endmodule



// megafunction wizard: %ALTPLL%
// ...
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
// ...

module pll ( inclk0, c0);

		input     inclk0;
        output    c0;

		wire [0:0] sub_wire2 = 1'h0;
        wire [4:0] sub_wire3;
        wire  sub_wire0 = inclk0;
        wire [1:0] sub_wire1 = {sub_wire2, sub_wire0};
        wire [0:0] sub_wire4 = sub_wire3[0:0];
        wire  c0 = sub_wire4;

        altpll altpll_component ( .inclk (sub_wire1), .clk
          (sub_wire3), .activeclock (), .areset (1'b0), .clkbad
          (), .clkena ({6{1'b1}}), .clkloss (), .clkswitch
          (1'b0), .configupdate (1'b0), .enable0 (), .enable1 (),
          .extclk (), .extclkena ({4{1'b1}}), .fbin (1'b1),
          .fbmimicbidir (), .fbout (), .fref (), .icdrclk (),
          .locked (), .pfdena (1'b1), .phasecounterselect
          ({4{1'b1}}), .phasedone (), .phasestep (1'b1),
          .phaseupdown (1'b1), .pllena (1'b1), .scanaclr (1'b0),
          .scanclk (1'b0), .scanclkena (1'b1), .scandata (1'b0),
          .scandataout (), .scandone (), .scanread (1'b0),
          .scanwrite (1'b0), .sclkout0 (), .sclkout1 (),
          .vcooverrange (), .vcounderrange ());

        defparam
                altpll_component.bandwidth_type = "AUTO",
                altpll_component.clk0_divide_by = 250,
                altpll_component.clk0_duty_cycle = 50,
                altpll_component.clk0_multiply_by = 1,
                altpll_component.clk0_phase_shift = "0",
                altpll_component.compensate_clock = "CLK0",
                altpll_component.inclk0_input_frequency = 20000,
                altpll_component.intended_device_family = "Cyclone IV E",
                altpll_component.lpm_hint = "CBX_MODULE_PREFIX=lab1clk",
                altpll_component.lpm_type = "altpll",
                altpll_component.operation_mode = "NORMAL",
                altpll_component.pll_type = "AUTO",
                altpll_component.port_activeclock = "PORT_UNUSED",
                altpll_component.port_areset = "PORT_UNUSED",
                altpll_component.port_clkbad0 = "PORT_UNUSED",
                altpll_component.port_clkbad1 = "PORT_UNUSED",
                altpll_component.port_clkloss = "PORT_UNUSED",
                altpll_component.port_clkswitch = "PORT_UNUSED",
                altpll_component.port_configupdate = "PORT_UNUSED",
                altpll_component.port_fbin = "PORT_UNUSED",
                altpll_component.port_inclk0 = "PORT_USED",
                altpll_component.port_inclk1 = "PORT_UNUSED",
                altpll_component.port_locked = "PORT_UNUSED",
                altpll_component.port_pfdena = "PORT_UNUSED",
                altpll_component.port_phasecounterselect = "PORT_UNUSED",
                altpll_component.port_phasedone = "PORT_UNUSED",
                altpll_component.port_phasestep = "PORT_UNUSED",
                altpll_component.port_phaseupdown = "PORT_UNUSED",
                altpll_component.port_pllena = "PORT_UNUSED",
                altpll_component.port_scanaclr = "PORT_UNUSED",
                altpll_component.port_scanclk = "PORT_UNUSED",
                altpll_component.port_scanclkena = "PORT_UNUSED",
                altpll_component.port_scandata = "PORT_UNUSED",
                altpll_component.port_scandataout = "PORT_UNUSED",
                altpll_component.port_scandone = "PORT_UNUSED",
                altpll_component.port_scanread = "PORT_UNUSED",
                altpll_component.port_scanwrite = "PORT_UNUSED",
                altpll_component.port_clk0 = "PORT_USED",
                altpll_component.port_clk1 = "PORT_UNUSED",
                altpll_component.port_clk2 = "PORT_UNUSED",
                altpll_component.port_clk3 = "PORT_UNUSED",
                altpll_component.port_clk4 = "PORT_UNUSED",
                altpll_component.port_clk5 = "PORT_UNUSED",
                altpll_component.port_clkena0 = "PORT_UNUSED",
                altpll_component.port_clkena1 = "PORT_UNUSED",
                altpll_component.port_clkena2 = "PORT_UNUSED",
                altpll_component.port_clkena3 = "PORT_UNUSED",
                altpll_component.port_clkena4 = "PORT_UNUSED",
                altpll_component.port_clkena5 = "PORT_UNUSED",
                altpll_component.port_extclk0 = "PORT_UNUSED",
                altpll_component.port_extclk1 = "PORT_UNUSED",
                altpll_component.port_extclk2 = "PORT_UNUSED",
                altpll_component.port_extclk3 = "PORT_UNUSED",
                altpll_component.width_clock = 5;


endmodule

